
`timescale 1ns/10ps
`celldefine
module TIEHL (tiehi, tielo);
output  tiehi ;
output  tielo ;

assign tiehi = 1'b1;
assign tielo = 1'b0;
endmodule
`endcelldefine

